module dadda_tree(
input [5:0]pp0, pp1, pp2, pp3, pp4, pp5, // 6 partial products
input [5:0]pp6, pp7, pp8, pp9, pp10, pp11, // 6 partial products
output 
);

endmodele